/*
 * Copyright © 2017-2020 Eric Matthews,  Lesley Shannon
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * Initial code developed under the supervision of Dr. Lesley Shannon,
 * Reconfigurable Computing Lab, Simon Fraser University.
 *
 * Author(s):
 *             Eric Matthews <ematthew@sfu.ca>
 */

package cva5_types;
    import cva5_config::*;
    import riscv_types::*;
    import csr_types::*;

    localparam FLEN_INTERNAL = 34;

    localparam LOG2_RETIRE_PORTS = $clog2(RETIRE_PORTS);
    localparam LOG2_MAX_IDS = $clog2(MAX_IDS);

    typedef logic[LOG2_MAX_IDS-1:0] id_t;
    typedef logic[1:0] branch_predictor_metadata_t;

    typedef logic [3:0] addr_hash_t;
    typedef logic [5:0] phys_addr_t;

    typedef struct packed {
        logic isFloat;
        rs_addr_t rs;
    } rf_addr_t;

    typedef enum logic [1:0] {
        ALU_CONSTANT = 2'b00,
        ALU_ADD_SUB = 2'b01,
        ALU_SLT = 2'b10,
        ALU_SHIFT = 2'b11
    } alu_op_t;

    typedef enum logic [1:0] {
        ALU_LOGIC_XOR = 2'b00,
        ALU_LOGIC_OR = 2'b01,
        ALU_LOGIC_AND = 2'b10,
        ALU_LOGIC_ADD = 2'b11
    } alu_logic_op_t;

    typedef struct packed{
        logic valid;
        exception_code_t code;
        logic [31:0] tval;
        logic [31:0] pc;
        id_t id;
    } exception_packet_t;

    typedef struct packed{
        logic ok;
        exception_code_t error_code;
    } fetch_metadata_t;

    typedef struct packed{
        id_t id;
        logic [31:0] pc;
        logic [31:0] instruction;
        logic valid;
        fetch_metadata_t fetch_metadata;
    } decode_packet_t;

    typedef struct packed{
        logic [31:0] pc;
        logic [31:0] instruction;
        logic [2:0] fn3;
        logic [6:0] opcode;

        rs_addr_t rd_addr;
        phys_addr_t phys_rd_addr;

        logic uses_rd;
        logic is_multicycle;
        id_t id;
        exception_sources_t exception_unit;
        logic stage_valid;
        fetch_metadata_t fetch_metadata;
    } issue_packet_t;

    typedef struct packed{
        logic [XLEN:0] in1;//contains sign padding bit for slt operation
        logic [XLEN:0] in2;//contains sign padding bit for slt operation
        logic [XLEN-1:0] shifter_in;
        logic [31:0] constant_adder;
        alu_op_t alu_op;
        alu_logic_op_t logic_op;
        logic [4:0] shift_amount;
        logic subtract;
        logic arith;//contains sign padding bit for arithmetic shift right operation
        logic lshift;
    } alu_inputs_t;

    typedef struct packed {
        logic [XLEN:0] rs1;
        logic [XLEN:0] rs2;
        logic [31:0] pc_p4;
        logic [2:0] fn3;
        logic [31:0] issue_pc;
        logic issue_pc_valid;
        logic jal;
        logic jalr;
        logic jal_jalr;
        logic is_call;
        logic is_return;
        logic [20:0] pc_offset;
    } branch_inputs_t;

    typedef struct packed {
        id_t id;
        logic valid;
        logic [31:0] pc;
        logic [31:0] target_pc;
        logic branch_taken;
        logic is_branch;
        logic is_return;
        logic is_call;
    } branch_results_t;

    typedef struct packed{
        logic [XLEN-1:0] rs1_load;
        logic [XLEN-1:0] rs2;
        logic [4:0] op;
    } amo_alu_inputs_t;

    typedef struct packed{
        logic is_lr;
        logic is_sc;
        logic is_amo;
        logic [4:0] op;
    } amo_details_t;

    typedef struct packed{
        logic [XLEN-1:0] rs1;
        logic [XLEN-1:0] rs2;
        logic [11:0] offset;
        logic [2:0] fn3;
        logic load;
        logic store;
        logic fence;
        logic forwarded_store;
        id_t store_forward_id;
        //amo support
        amo_details_t amo;
    } load_store_inputs_t;

    typedef struct packed{
        logic [XLEN-1:0] rs1;
        logic [XLEN-1:0] rs2;
        logic [1:0] op;
    } mul_inputs_t;

    typedef struct packed{
        logic [XLEN-1:0] rs1;
        logic [XLEN-1:0] rs2;
        logic [1:0] op;
        logic reuse_result;
    } div_inputs_t;

    typedef struct packed{
        csr_addr_t addr;
        logic[1:0] op;
        logic reads;
        logic writes;
        logic [XLEN-1:0] data;
    } csr_inputs_t;

    typedef enum logic [2:0] { 
        ORG_A_SIGN = 3'b000,
        ORG_B_SIGN = 3'b001,
        INV_A_SIGN = 3'b010,
        INV_B_SIGN = 3'b011,
        XOR_SIGNS = 3'b100
    } sign_mod_t;

    typedef struct packed { // -?((rs1(*rs2)?)|rs1) (+ -?(rs3|rs2))?
        logic mul; // rs1 * rs2. Result if none of the add-options is set
        logic add_mul_rs3; // result is (res of mul) + rs3
        logic add_rs1_rs2; // result rs1 + rs2
        sign_mod_t ovr_1st_add_in_sign; // changes sign bit of first add operand or result if none of the above result-modes is active
        logic negate_2nd_add_in; // flips sign bit of second add operand
    } fpmac_op_t;

    typedef enum logic [2:0] {
        FPMAC_OP = 3'b000,
        FPDIV_OP = 3'b001,
        FPSQRT_OP = 3'b010,
        FP_FROM_IEEE_OP = 3'b011,
        FPCVT_FROM_I_OP = 3'b100,
        FPCVT_FROM_U_OP = 3'b101,
        FPMIN_OP = 3'b110,
        FPMAX_OP = 3'b111
    } fpu_op_t;

    typedef struct packed{
        logic [FLEN_INTERNAL-1:0] rs1;
        logic [XLEN-1:0] rs1_gp;
        logic [FLEN_INTERNAL-1:0] rs2;
        logic [FLEN_INTERNAL-1:0] rs3;
        fpmac_op_t fpmac_op;
        fpu_op_t op;
    } fpu_inputs_t;

    typedef enum logic [2:0] {
        FP_TO_IEEE_OP = 3'b000,
        FPCVT_TO_I_OP = 3'b010,
        FPCVT_TO_U_OP = 3'b011,
        FPEQ_OP = 3'b100,
        FPLT_OP = 3'b101,
        FPLE_OP = 3'b110,
        FPCLASS_OP = 3'b111
    } fp_to_gp_op_t;

    typedef struct packed{
        logic [FLEN_INTERNAL-1:0] rs1;
        logic [FLEN_INTERNAL-1:0] rs2;
        fp_to_gp_op_t op;
    } fp_to_gp_inputs_t;

    typedef struct packed{
        logic [31:0] pc_p4;
        logic is_ifence;
        logic is_mret;
        logic is_sret;
    } gc_inputs_t;

    typedef struct packed {
        logic [31:0] addr;
        logic load;
        logic store;
        logic [3:0] be;
        logic [2:0] fn3;
        logic [31:0] data;
        id_t id;
        logic forwarded_store;
        id_t id_needed;
    } lsq_entry_t;

    typedef struct packed {
        logic [31:0] addr;
        logic [3:0] be;
        logic [2:0] fn3;
        logic forwarded_store;
        logic [31:0] data;
    } sq_entry_t;

    typedef struct packed {
        logic sq_empty;
        logic no_released_stores_pending;
        logic idle;
    } load_store_status_t;

    typedef struct packed{
        id_t id;
        logic valid;
        logic [MAX_POSSIBLE_REG_BITS-1:0] data;
    } wb_packet_t;

    typedef struct packed{
        id_t id;
        logic valid;
        phys_addr_t phys_addr;
        logic [MAX_POSSIBLE_REG_BITS-1:0] data;
    } commit_packet_t;

    typedef struct packed{
        logic valid;
        id_t phys_id;
        logic [LOG2_RETIRE_PORTS : 0] count;
    } retire_packet_t;

    typedef struct packed {
        logic [31:0] addr;
        logic load;
        logic store;
        logic [3:0] be;
        logic [2:0] fn3;
        logic [31:0] data_in;
        id_t id;
    } data_access_shared_inputs_t;

    typedef enum  {
        LUTRAM_FIFO,
        NON_MUXED_INPUT_FIFO,
        NON_MUXED_OUTPUT_FIFO
    } fifo_type_t;

    typedef struct packed{
        logic init_clear;
        logic fetch_hold;
        logic issue_hold;
        logic fetch_flush;
        logic writeback_supress;
        logic retire_hold;
        logic sq_flush;
        logic tlb_flush;
        logic exception_pending;
        exception_packet_t exception;
        logic pc_override;
        logic [31:0] pc;
    } gc_outputs_t;

    typedef struct packed {
        logic software;
        logic timer;
        logic external;
    } interrupt_t;
    
    typedef struct packed {
        //Fetch
        logic early_branch_correction;

        //Decode
        logic operand_stall;
        logic unit_stall;
        logic no_id_stall;
        logic no_instruction_stall;
        logic other_stall;
        logic instruction_issued_dec;
        logic branch_operand_stall;
        logic alu_operand_stall;
        logic ls_operand_stall;
        logic div_operand_stall;

        // Instruction mix
        logic alu_op;
        logic branch_or_jump_op;
        logic load_op;
        logic store_op;
        logic mul_op;
        logic div_op;
        logic misc_op;
        logic float_op;

        // Branch Prediction
        logic branch_correct;
        logic branch_misspredict;
        logic return_correct;
        logic return_misspredict;

        //Load Store Unit
        logic load_conflict_delay;
        logic ls_is_peri_access;

        //Register File
        logic rs1_forwarding_needed;
        logic rs2_forwarding_needed;
        logic rs1_and_rs2_forwarding_needed;

        // Instr. Invalidation
        logic instr_inv_stall;

        // Branch Results/Effects
		logic br_branch_taken;
		logic br_is_branch;
		logic br_is_return;
		logic br_is_call;
    } cva5_trace_events_t;

    typedef struct packed {
        logic [31:0] pc;
        logic [31:0] instruction;
        logic valid;
    } trace_retire_outputs_t;

    typedef struct packed {
        logic [31:0] instruction_pc_dec;
        logic [31:0] instruction_data_dec;
        logic [1:0] current_privilege;
        logic [31:0] branch_target_pc;
        cva5_trace_events_t events;
    } trace_outputs_t;


    typedef enum logic [11:0] {
        MINSTR_INV_CSR = 12'h7C0
    } cva5_csr_reg_addr_t;

endpackage
